module pulses; // Incorrect pulse generation attempt
  reg [8:0] I;
  reg a,b;