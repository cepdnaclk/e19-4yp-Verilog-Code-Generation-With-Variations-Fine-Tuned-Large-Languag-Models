module and