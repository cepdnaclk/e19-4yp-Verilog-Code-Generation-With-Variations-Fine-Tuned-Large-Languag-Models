module tst_dff_p_b();
  reg di,clk; wire do;
  dff_p d1(do,di,clk); //