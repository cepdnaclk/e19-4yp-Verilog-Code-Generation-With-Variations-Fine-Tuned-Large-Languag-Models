module AndOr (output X, Y, input A, B, C);
bit [7:0] A;
bit [7:0] B;
bit [7:0] C;
bit X;
bit Y;