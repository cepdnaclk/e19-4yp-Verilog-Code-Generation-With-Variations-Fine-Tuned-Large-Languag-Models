module tst_wand2_v; //testbench
reg i1,i2;
wire o; // Added wire declaration
wand2 ww(i1,i2,o);
initial
begin
i1=0; i2=0; // Drv1=pull0, Drv2=pull0 -> o = pull0 (wand rule)
end
initial $monitor($time,"i1=%b,i2=%b,o=%b",i1,i2,o);