module enum_strength (a, c, zn, zp);
input a, c;
output [1:0] zn, zp;
nmos (zn, a,