module Problem3();
output [3:0] out;
reg [3:0] A;
reg [3:0] B