module Ripple_Add;
    parameter COUNTER_WIDTH = 3;
    parameter ARRAY_LENGTH =