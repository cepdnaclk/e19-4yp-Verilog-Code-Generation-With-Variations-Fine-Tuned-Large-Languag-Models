module reg4(D, Clock, Resetn, Q);
input [3:0] D;
input Clock, Resetn;
output [3:0] Q;
reg [3:0] Q;
always @(posedge Clock or negedge Resetn)
    if (Resetn == 0)
        Q <= 4'b0000;
    else
        Q <= D;
endmodule
```

#### Cause

An array variable is declared inside an `if-else` conditional statement, and the `size` of the array is not specified.

#### Resolution

An array element must be accessed through a constant index, or an index value must be assigned to a variable.

#### References

* [IEEE P16