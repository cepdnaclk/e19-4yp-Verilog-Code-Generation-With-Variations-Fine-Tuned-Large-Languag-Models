`timescale 1ns/100ps
module ALU8 (input [7:0] left, right, input [1:0] mode, output reg [7:0] ALUout);
always_comb begin
    case (mode)
        0: ALUout = left + right;
        1: ALUout = left - right;
        2: ALUout = left & right;
        3: ALUout = left | right;
        default: ALUout = 8'bX;
    endcase
end
endmodule
### RTL Code:
![RTL code](https://github.com/Ayush8111/FINAL_PROJECT/blob/main/ALU_8bit_RISCV/RTL%20code.png)

### Coverage:
![Coverage](https://github.com/Ayush8111/FINAL_PROJECT/blob/main/ALU_8bit_RISCV/Coverage.png)
### Synthesis:
![Synthesis](https://github.com/Ayush8111/FINAL_PROJECT/blob/main/ALU_8bit_RISCV/synth.PNG)
### RTL Code:
![RTL Codes](https://github.com/Ayush8111/FINAL_PROJECT/blob/main/ALU_8bit_RISCV/RTL%