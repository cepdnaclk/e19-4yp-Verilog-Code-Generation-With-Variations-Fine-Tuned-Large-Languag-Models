module latch_