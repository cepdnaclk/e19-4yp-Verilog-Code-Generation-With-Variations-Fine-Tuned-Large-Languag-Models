module g(a,a1,b,c,b1,c1);
input b,c,b1,c1;
output [15:0] a;
wire [15:0] a1;
wire [15:0]