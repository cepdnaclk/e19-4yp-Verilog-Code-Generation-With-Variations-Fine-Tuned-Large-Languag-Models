module Problem1(input [3:0] a, b, output [3:0] sum);
  logic di, clk;
  integer x, y, sum;