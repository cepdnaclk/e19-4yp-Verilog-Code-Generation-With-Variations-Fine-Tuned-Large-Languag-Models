module AndOr (output X, Y, input A, B, C);
`ifdef USE_BIT_INPUT
bit A, B, C;
`else
wire A, B, C;
`endif
assign #10 X = A & B;
assign #10 Y = B | C;
endmodule
### Result:
#### Run with USE_BIT_INPUT defined
+------+----------------------+----------------------+
| Name | Original Module      | Modified Module      |
+------+----------------------+----------------------+
| A    | 0                    | 0                    |
+------+----------------------+----------------------+
| B    | 0                    | 0                    |
+------+----------------------+----------------------+
| C    | 0                    | 0                    |
+------+----------------------+----------------------+
| X    | 0                    | 0                    |
+------+----------------------+----------------------+
| Y    | 0                    | 0                    |
+------+----------------------+----------------------+
#### Run with USE_BIT_INPUT not defined
+------+----------------------+---------------------+
| Name | Original Module      | Modified Module     |
+------+----------------------+---------------------+
| A    | 0                    | 0                   |
+------+----------------------+---------------------+
| B    | 0                    | 0                   |
+------+----------------------+---------------------+
| C    | 0                    | 0                   |
+------+----------------------+---------------------+
| X    | 0                    | 0                   |
+------+----------------------+---------------------+
| Y    | 0                    | 0                   |
+------+----------------------+---------------------+
### Version Requirement
| OCaml version | Opam package version |
|--------------|----------------------|