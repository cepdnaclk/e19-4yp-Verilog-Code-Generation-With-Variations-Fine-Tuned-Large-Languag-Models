```
module aoi3_2(g1,g2,a,b,c