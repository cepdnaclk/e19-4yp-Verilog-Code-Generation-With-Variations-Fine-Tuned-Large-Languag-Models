module tst_CMOSsw1();
  reg in,con; wire out;
  CMOSsw1 cmsw[2:0](out[1:0],in,con); // Instantiate CMOS switch
  initial begin in=1'b0; con=1'b1; end // Start enabled
  always #5 in =~in; // Toggle data
  always #3 con=~con; // Toggle control
  initial $monitor($time, "in = %b, con = %b, output = %b ",in,con,out);
  initial #20 $stop; // Stop simulation
  initial
  begin
    for(i=0;i<3;i=i+1)
    begin
        $display("in = %b, con = %b, output = %b ",in,con,out