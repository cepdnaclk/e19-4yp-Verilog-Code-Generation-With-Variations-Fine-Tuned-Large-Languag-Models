timescale 1ns/100ps
module maj3 (
    input a, b, c, output y
);
wire im1, im2, im3;
parameter
    tplh1=2, tphl1=4