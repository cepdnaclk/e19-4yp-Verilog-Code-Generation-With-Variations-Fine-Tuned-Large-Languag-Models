module dff(do,di,clk); // Behavioral D Flip-Flop
output [3:0] do;
input [3:0] di