module ror (d, clock, input);
input [3:0] d, clock