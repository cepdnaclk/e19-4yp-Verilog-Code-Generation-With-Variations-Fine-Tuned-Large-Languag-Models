module wire_assign( input in, output logic out );
    // assign out to in
    assign out = in;
endmodule
### Result:
The new code should pass simulations.