module IR_DV (input logic [7:0] data_in, input logic load, clk,
output reg [7:0] data_out);
// Create a 7