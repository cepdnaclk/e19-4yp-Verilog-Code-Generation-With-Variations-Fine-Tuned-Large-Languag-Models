module full_adder(i1, i2, cin, sum, cout);
input i1, i2, cin;
output [1:0] sum, cout;
assign sum =