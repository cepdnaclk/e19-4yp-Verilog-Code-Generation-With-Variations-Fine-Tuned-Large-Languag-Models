module gade(a,a1,b,c,b1,c1);
input b