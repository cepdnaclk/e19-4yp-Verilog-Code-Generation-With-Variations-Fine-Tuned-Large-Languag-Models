module Problem10(input [3:0] a, b