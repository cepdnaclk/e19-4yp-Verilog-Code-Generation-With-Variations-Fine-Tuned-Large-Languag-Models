module pulses