module testbench ();
data a = {
    x: rand
};
generate a;
process a