module tstha_10(clk,rst,a,b,ca,s);