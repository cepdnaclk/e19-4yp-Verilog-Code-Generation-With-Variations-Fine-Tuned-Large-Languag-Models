module example6(x1, x2, x3, x4, f, g, h);
input x1, x2, x3, x4;