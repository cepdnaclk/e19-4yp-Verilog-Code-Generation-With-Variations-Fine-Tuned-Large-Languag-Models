module AndOr (output X, Y, input A, B, C);
wire