module testbench ();
generate struct begin