```verilog
module tst_mup; // Testbench for Microprocessor
reg clk,en,int; // Clock, Enable, Interrupt inputs
// Assuming mup_opr is the microprocessor module instance
mup_opr rr(clk,int,en); // Instantiate DUT
initial
begin
int=1'b0;clk=1'b0;en=1'b0; // Initialize
end
always #2 clk=~clk; // Generate clock
// Monitor clock, time, inputs, and internal MUP registers (pc, ir, dcop)
initial $monitor("clk=%b, t=%0d, en=%b, int=%b, rr.pc=%0d, rr.ir=%0h, rr.dcop=%0d", clk,$time,en,int,rr.pc,rr.ir,rr.dcop); // Corrected format specifiers
// mup_opr rr(clk,int,en); // Instantiate DUT
initial #40 $stop; // Stop simulation
endmodule
```
### Result of Testing:
#### Corrected `pkg::consts[BCD_in]`:
![Corrected `pkg::consts[BCD_in]`](https://github.com/DengyuanZ