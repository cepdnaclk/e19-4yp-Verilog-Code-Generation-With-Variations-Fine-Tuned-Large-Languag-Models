module test;
wire [31:0] a[0:7];
wire [31:0] b[0:7];
wire [31:0] c[0:7];
wire [31:0] d[0:7];
wire [31:0] e[0:7];
wire [31:0] f[0:7];
wire [31:0] g[0:7];
wire [31:0] h[0:7];
wire [31:0] i[0:7];
wire [31:0] j[0:7];
wire [31:0] k[0:7];
wire [31:0] l[0:7];
wire [31:0] m[0:7];
wire [31:0] n[0:7];
wire [31:0] o[0:7];
wire [31:0] p[0:7];
wire [31:0] q[0:7];
wire [31:0] r[0:7];
wire [31:0] s[0:7];
wire [31:0] t[0:7];
wire [31:0] u[0:7];
wire [31:0] v[0:7];
wire [31:0] w[0:7];
wire [31:0] x[0:7];
wire [31:0] y[0:7];
wire [31:0] z;
initial begin
    a[0] = 1'b0;
    a[1] = 1'b1;
    a[2] = 1'b0;
    a[3] = 1'b1;
    a[4] = 1'b0;
    a[5] = 1'b0;
    a[6] = 1'b1;
    a[7] = 1'b1;
    b[0] = 1'b0;
    b[1] = 1'b1;
    b[2] = 1'b0;
    b[3] = 1'b1;
    b[4] = 1'b0;
    b[5] = 1'b0;
    b[6] = 1'b1;
    b[7] = 1'b1;
    c[0] = 1'b0;
    c[1] = 1'b1;
    c[2] = 1'b1;
    c[3] = 1'b0;
    c[4] = 1'b0;
    c[5] = 1'b0;
    c[6] = 1'b1;
    c[7] = 1'b1;
end
always @*
    d[0] = a[0] ^ a[1] ^ a[4];
    d[1] = a[1] ^ a[2] ^ a[5];
    d[2] = a[2] ^ a[3] ^ a[6];
    d[3] = a[3] ^ a[4] ^ a[7];
    d[4] = a[4] ^ a[5] ^ a[0];
    d[5] = a[5] ^ a[6] ^ a[1];
    d[6] = a[6] ^ a[7] ^ a[2];
    d[7] = a[7] ^ a[0] ^ a[3];
    e[0] = a[0] & a[1] & a[4];
    e[1] = a[1] & a[2] & a[5];
    e[2] = a[2] & a[3] & a[6];
    e[3] = a[3] & a[4] & a[7];
    e[4] = a[4] & a[5] & a[0];
    e[5] = a[5] & a[6] & a[1];
    e[6] = a[6] & a[7] & a[2];
    e[7] = a[7] & a[0] & a[3];
    f[