module EventCtlPart (output xPart, yPart, input a, b, c);
reg xReg, yReg;
assign xPart = xReg;
assign yPart = yReg;
always @(a, b)
begin: PartList
    xReg <= a & b & c;
    if (b) begin
        if (c) begin
            yReg <= 1'b1;
        end
        else begin
            yReg <= 1'b0;
        end
    end
    else