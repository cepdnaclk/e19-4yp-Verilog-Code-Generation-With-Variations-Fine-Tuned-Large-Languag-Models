module TOP1 (CLK, RST_X, OUTP);

  input CLK, RST_X;
  output OUTP;
  wire [7:0] inp0 = 8'h50;
  wire [7:0] inp1 = 8'h60;

  wire [7:0] x;
  wire [7:0] y;

  always @ (posedge CLK) begin
    x <= RST_X? 8'h10 : x + 1;
    y <= RST_X? 8'h20 : y + 1;
  end

  wire outp;
  assign outp = inp0 inside {8'h10, 8'h20, 8'h30};

  assign OUTP = outp;
endmodule
### Modified Top Module Instantiation:
module tb_TOP1;
  reg CLK, RST_X;
  TOP1 uut(.CLK(CLK),.RST_X(RST_X));
  initial begin
    CLK = 0;
    forever #5 CLK = ~CLK;
  end

  initial begin
    RST_X = 0; #10;
    RST_X = 1;
  end
endmodule
### Modified Package:
package com_p;
    parameter COMPARE_W = 8;
    parameter COMPARE_L = 3;
    constant comparators [COMPARE_L-1:0][COMPARE_W-1:0] = {8'h10, 8'h20, 8'h30};
endpackage
### Expected Output:
### -----------------------------
### Output #1 (for `outp` = 1):
### -----------------------------
*X*
### -----------------------------
### Output #2 (for `outp` = 0):
### -----------------------------
X
### -----------------------------
### Output #3 (for `outp` = 0):
### -----------------------------
X
### -----------------------------
### Output #4 (for `outp` = 0):
### -----------------------------
X
### -----------------------------
### Output #5 (for `outp` = 0):
### -----------------------------
X
### -----------------------------
### Output #6 (for `outp` = 0):
### -----------------------------
X
### -----------------------------
### Output #7 (for `outp` = 0):
### -----------------------------
X
### -----------------------------
### Output #8 (for `outp` = 0):
### -----------------------------
X
### -----------------------------
### Output #9 (for `outp` = 0):
### -----------------------------
X
### -----------------------------
### Output #10 (for `outp` = 0):
### -----------------------------
X
### -----------------------------
### Output #11 (for `outp` = 0):
### -----------------------------
X
### -----------------------------
### Output #12 (for `outp` = 0):
### -----------------------------
X
### -----------------------------
### Output #13 (for `outp` = 0):
### -----------------------------
X
### -----------------------------
### Output #14 (for `outp` = 0):
### -----------------------------
X
### -----------------------------
### Output #15 (for `outp` = 0):
### -----------------------------
X
### -----------------------------
### Output #16 (for `outp` = 0):
### -----------------------------
X
### -----------------------------
### Output #17 (for `outp` = 0):
### -----------------------------
X
### -----------------------------
### Output #18 (for `outp` = 0):
### -----------------------------
X
### -----------------------------
### Output #19 (for `outp` = 0):
### -----------------------------
X
### -----------------------------
### Output #20 (for `outp` = 0):
###