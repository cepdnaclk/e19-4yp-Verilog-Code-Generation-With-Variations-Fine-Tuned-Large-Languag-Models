module gade(a,a1,b,c,b1,c1);
input b,c,b1,c1;
output [2:0] a,a1;
// Instantiate OR gate with inertial delay 3
or #3 gg1(a1[2],c1,b1);
// Instantiate AND gate with rise=2, fall=1 inertial delay
and #(2,1) gg2(a[1:0],c,b);
endmodule
module gade(a,a1,b,c,b1,c1);
input b,c,b1,c1;
output [2:0] a,a1;
// Instantiate OR gate with inertial delay 3
or #3 gg1(a1[2],c1,b1);
// Instantiate AND gate with rise=2, fall=1 inertial delay
and #(2,1) gg2(a[1:0],c,b);
endmodule

### Base Verilog