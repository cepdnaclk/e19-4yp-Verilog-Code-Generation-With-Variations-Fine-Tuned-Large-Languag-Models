module tstha_10();
  reg a,