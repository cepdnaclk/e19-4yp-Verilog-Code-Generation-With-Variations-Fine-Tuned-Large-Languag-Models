module tstha_9();
  reg [3:0] clk; wire s,ca;