```verilog
// Create the module
module reg