module RAM4 (output[7:0] Obus, input[7:0] Ibus, input[3:0] Ad