module tst