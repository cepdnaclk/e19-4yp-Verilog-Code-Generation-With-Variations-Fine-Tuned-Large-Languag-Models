module example9(x1, x2, x3, f);
input x1, x2, x3;
output f;
reg f;
always @(x1 or