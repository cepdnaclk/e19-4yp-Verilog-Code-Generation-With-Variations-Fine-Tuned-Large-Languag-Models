module ha_4(s,ca,a,b); // Half Adder with gate delays
  input