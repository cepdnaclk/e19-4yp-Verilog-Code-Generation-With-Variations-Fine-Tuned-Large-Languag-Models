module tst_alu4();
  reg [3:0]a,b; reg[1:0] f; reg cci; wire[3:0]d