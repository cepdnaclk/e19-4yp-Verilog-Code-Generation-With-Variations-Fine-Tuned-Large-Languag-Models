module gade(a,a1,b,c,b1,c1);
input b,c,b1,c1;
output a,a1;
// Instantiate OR gate with inertial delay 3
or #3 gg1(a1,c1,b1);
// Instantiate AND gate with rise=2, fall=1 inertial delay
and #(2,1) gg2(a,c,b);
endmodule
### Compilation
`ncvlog gade.v`
### Running Simulation
##### Output:
`ncvlog: *E,UNHANDLED (Unhandled statement)`
`ncvlog: *W,NCEG2003 (Naming Conventions: Inconsistent naming between `gade.v' and unnamed item in file: