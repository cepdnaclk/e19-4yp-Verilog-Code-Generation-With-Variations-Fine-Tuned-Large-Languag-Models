module AndOr (output