module Ripple_Add;
    FA fa0();