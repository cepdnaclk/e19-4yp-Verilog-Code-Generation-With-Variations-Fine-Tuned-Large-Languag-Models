module gates4 (
input wire [3:0] x,
output wire [3:0]