module display(in, out);
struct packed {
logic [7:0] in;
logic out