module aoi_gate(o,a1,a2,b1,b2);
input a1,a2,b1,b2;// a1,a2,b1,b2 form the input
//ports of the module
output [3:0] o;//o is the single output port of the module
wire [3:0] o1,o2;//o1 and o2 are intermediate signals
//within the module
and g1(o1,a1,a2); //The AND gate primitive has two
and g2(o2,b1,b2);// instantiations with assigned
//names g1 & g2.
nor g3(o[0],o1,o2);//The nor gate has one instantiation
//with assigned name g3.
endmodule

### Output File: