module example_module;
  logic [3:0]