module DataComponent (DataIn, DataOut, ControlSignals);
input [7:0] Data