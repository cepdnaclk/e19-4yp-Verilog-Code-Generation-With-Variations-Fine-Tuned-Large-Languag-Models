module tst_up