module example3(Data, Clock, Reset, RegSum, Sum);
input Clock, Reset;
input [3:0