module counter (
     input wire cl