module test(dout,din