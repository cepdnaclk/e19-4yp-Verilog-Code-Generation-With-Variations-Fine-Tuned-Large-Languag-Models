module par(in, parity, all_ones);
  struct {
    logic [7:0] x1;
    logic [7:0] x2;
    logic [7:0] x3;
    logic [7:0] x4