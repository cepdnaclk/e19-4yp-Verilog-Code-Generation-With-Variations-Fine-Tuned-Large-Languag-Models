module wire_assign( input bit in, output out );
    // assign out to in
    assign out = in;
endmodule
### Result of Test
Test Passed
*/



module wire_assign( input bit in, output out );
    // assign out to in
    assign out = in;
endmodule