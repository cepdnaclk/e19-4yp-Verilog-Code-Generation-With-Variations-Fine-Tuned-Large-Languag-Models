module aoibeh2(o,a,b); // Mixed structural/behavioral AOI
output o;
input[1:0]a,b;
wire a1,b1; // Outputs of AND gates
reg o; // Behavioral output must be reg
// Structural AND gates using primitives
and g1(a1,a[1],a[0]), g2(b1,b[1],b[0]);
// Behavioral NOR logic sensitive to AND outputs
always@(a1 or b1)
o = ~(a1 || b1);
initial begin : foo
  o <= {4{1'b0}};
  o[0] <= 1'b1;
  #10;
  o[1] <= 1'b1;
  #10;
  #30;
  o[2] <= 1'b1;
  #10;
  #30;
  o[3] <= 1'b1;
  #10;
  #30;
  #100;
  o[1] <= 1'b0;
  #30;
  #100;
  o[1] <= 1'b1;
  #50;
  o[0] <= 1'b0;
  #30;
  #100;
  o[0] <= 1'b1;
  #50;
  o[1] <= 1'b0;
  #50;
  o[2] <= 1'b0;
  #50;
  o[3] <= 1'b0;
  #100;
  #200;
  o[0] <= 1'b1;
  #50;
  o[1] <= 1'b1;
  #100;
  #200;
  o[0] <= 1'b0;
  #200;
  #200;
  o[1] <= 1'b0;
  #200;
  o[0] <= 1'b1;
  #200;
  o[1] <= 1'b1;
  #200;
  o[3] <= 1'b1;
  #200;
  #200;
  o[3] <= 1'b0;
  #200;
  o[2] <= 1'b1;
  #200;
  o[3] <= 1'b1;
  #200;
  o[2] <= 1'b0;
  #200;
  o[0] <= 1'b0;
  #200;
  o[1] <= 1'b0;
  #200;
  o[0] <= 1'b1;
  #200;
  o[0] <= 1'b0;
  #200;
  o[1] <= 1'b1;
  #200;
  o[1] <= 1'b0;
  #200;
  o[2] <= 1'b1;
  #200;
  o[1] <= 1'b1;
  #200;
  o[1] <= 1'b0;
  #200;
  o[3] <= 1'b1;
  #200;
  o[3] <= 1'b0;
  #200;
  o[2] <= 1'b1;
  #200;
  o[0] <= 1'b1;
  #200;
  o[1] <= 1'b0;
  #200;
  o[0] <= 1'b0;
  #200;
  o[2] <= 1'b1;
  #200;
  o[3] <= 1'b1;
  #200;
  o[3] <= 1'b0;
  #200;
  #900;
end : foo
end