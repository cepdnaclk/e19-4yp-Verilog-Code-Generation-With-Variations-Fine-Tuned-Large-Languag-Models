module gates4_top (
input wire [3:0] sw,
output wire [2:0] ld
);
wire