module contres(o,i1,i2);
input i1,i2;
output o;
// Drive wire 'o' from two buffers with