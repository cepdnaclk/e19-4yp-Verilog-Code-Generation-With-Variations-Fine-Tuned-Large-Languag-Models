module example7_10(x1, x2, x3, Clock, f, g);
input x1, x2, x3, Clock;
output f, g;