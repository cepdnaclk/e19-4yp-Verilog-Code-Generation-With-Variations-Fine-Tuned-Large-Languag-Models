module tst_wand1; //testbench
reg i1,i