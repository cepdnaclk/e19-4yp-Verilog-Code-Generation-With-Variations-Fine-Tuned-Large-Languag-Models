module test;
wire a;
wire [3:0] x;
wire [3:0] y;
wire [3:0] z;
struct {
    logic x