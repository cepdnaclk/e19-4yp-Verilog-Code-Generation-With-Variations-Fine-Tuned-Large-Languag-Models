module ripple_carry_1(cin,x,