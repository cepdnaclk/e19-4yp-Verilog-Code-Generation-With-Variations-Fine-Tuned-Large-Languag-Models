module func2(x