module for_if(i); logic i;
// A for loop with a if condition
// Nested in an if block to break out of the for loop
if (1) begin
    for (i = 0; i < 3; i = i