module example7_5mod3(x1, x2, x3