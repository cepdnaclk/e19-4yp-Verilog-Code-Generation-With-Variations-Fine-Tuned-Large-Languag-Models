module wire_assign( input in, output out );
    reg f;
    // assign out to in
    assign out = in