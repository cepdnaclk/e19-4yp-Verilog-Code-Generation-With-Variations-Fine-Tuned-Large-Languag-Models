module aoibeh2_6(o,a,b); // AOI w/ intial block
output o;
input[1:0]a,b;
wire a1,b1; // Outputs of AND gates