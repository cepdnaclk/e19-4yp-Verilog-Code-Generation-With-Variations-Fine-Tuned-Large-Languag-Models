module Problem8tb();
  Problem8 dut(.a(a),.b(b),