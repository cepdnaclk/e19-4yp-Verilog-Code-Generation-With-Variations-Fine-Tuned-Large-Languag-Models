module tst_wand7; //testbench
reg i1[7:0],i2[7:0];
wire