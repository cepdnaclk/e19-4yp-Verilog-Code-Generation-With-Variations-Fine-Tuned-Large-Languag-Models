module clock_gen_for_loop; // Renamed module for clarity
  reg clk, en;