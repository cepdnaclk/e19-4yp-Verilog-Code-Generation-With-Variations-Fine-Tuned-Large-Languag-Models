module tb_dff();
logic CLK, RESETn;
logic D, Q;
integer index;
logic [7:0] test_vectors