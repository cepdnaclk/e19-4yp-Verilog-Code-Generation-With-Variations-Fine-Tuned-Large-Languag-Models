module latch (input d