module ALU ( input [7:0] a, b, input pass, add,