module tst_ctr