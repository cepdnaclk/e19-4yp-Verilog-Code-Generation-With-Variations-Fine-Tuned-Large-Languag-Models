module test_enum (a,b,c,d,e,f,g,h,i,j,k,l,m,n);
	parameter x = 3, y = 3, z = 1;
	output a,b,c,d,e,f,g,h,i,j,k,l,m,n;
	input [2:0] c,d,e,f,g,h,i,j,k,l,m,n;
	wire abcd = a && b && c && d;
	wire abce = a && b && c && e;
	wire abcf = a && b && c && f;
	wire abcg = a && b && c && g;
	wire abch = a && b && c && h;
	wire abci = a && b && c && i;
	wire abcj = a && b && c && j;
	wire abcj = a && b && c && k;
	wire abcj = a && b && c && l;
	wire abcj = a && b && c && m;
	wire abcj = a && b && c && n;
	wire abcd = a && b && d;
	wire abce = a && b && e;
	wire abcf = a && b && f;
	wire abcg = a && b && g;
	wire abch = a && b && h;
	wire abci = a && b && i;
	wire abcj = a && b && j;
	wire abcj = a && b && k;
	wire abcj = a && b && l;
	wire abcj = a && b && m;
	wire abcj = a && b && n;
	wire abcd = a && b && c;
	wire abce = a && b && d;
	wire abcf = a && b && e;
	wire abcg = a && b && f;
	wire abch = a && b && g;
	wire abci = a && b && h;
	wire abcj = a && b && i;
	wire abcj = a && b && j;
	wire abcj = a && b && k;