module latch (input d, c, output reg q, q_b );