module tst_alu1();
  reg [3:0]a,b; reg[3:0] c; reg[2:0] f; reg cci; wire[3:0]d; wire co;
  alu_1 aa(d,co,a,b,f,