module testbench ();
    struct {
        logic [3:0] rand;
    } data;
generate data;
process data;
endmodule
### Expected Output:
```