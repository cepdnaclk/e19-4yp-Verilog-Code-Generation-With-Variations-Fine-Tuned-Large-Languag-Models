reg [