module DFF (input logic clk, rst, input logic [1:0] din, output logic [