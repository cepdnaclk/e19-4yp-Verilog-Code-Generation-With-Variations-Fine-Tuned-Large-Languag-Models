module AndOr (output X, Y, input A, B, C);
assign X = A & B;
assign Y = B | C;
end