module example4(x1, x2, x3, x4, f, g, h);