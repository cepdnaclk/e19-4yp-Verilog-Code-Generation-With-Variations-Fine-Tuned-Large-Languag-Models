```
module or_gate(b,a,en);
parameter N = 4;
input [N-1:0] a;
input en