module tst_alu4();
  reg [3:0]a,b; reg[1:0] f; reg cci; logic[3:0]d; logic co;
  //alu_4 aa(d,co,a,b,f,cci);
  always_comb begin // Instantiate ALU
  end
  initial $monitor($time, " cci = %b, a= %h,b = %