module SchedDelayL;
reg a, b;
initial
begin
end
always @(b) a = b