module test;
struct packed {
    logic x;