Modify the code at line 19 to line 33 to include a 4-bit data width. The code must generate a 4-bit long shift register.
```
module dff_4_inst(D, Clock, Resetn, Q);
input [3:0] D;
input Clock;
input Resetn;
output [3:0] Q;
integer i;
integer N;
initial N = 4;
reg [3:0] Q_reg;
always @