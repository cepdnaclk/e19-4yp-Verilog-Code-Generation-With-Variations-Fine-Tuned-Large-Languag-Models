`timescale 1ns/100ps
module maj4 (input [2:0] a, output reg [1