module test;
wire a;
union {logic x, y, z;} x