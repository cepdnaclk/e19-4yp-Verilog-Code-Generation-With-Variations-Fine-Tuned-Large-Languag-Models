```cpp
module AndOr (output X, Y, input [1:0] A, B, C);
assign #1