module ALU (input[3:0] ArgA, ArgB, input Clk, output logic Result, input Clock);
specify
    specparam tRise =