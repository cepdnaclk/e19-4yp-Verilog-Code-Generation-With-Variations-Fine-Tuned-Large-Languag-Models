module jk(clk,rst,set,d,q);
  input clk,rst,set,d;
  output q;
  reg q;