`timescale 1ns/100ps

module ShiftRegister32 (input sl, sr