module netdelay2(x,y);
input x;