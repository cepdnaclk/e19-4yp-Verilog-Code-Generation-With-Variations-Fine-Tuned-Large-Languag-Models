module tst_dff_p_b();
  reg di,clk; wire do;
  dff_p d1[2](do,di,clk); // Instantiate the DFF
  initial begin clk=0; di=1'b0; #35 $stop; end // Initialize & stop
  always #3 clk=~clk; // Generate clock
  always #5 di=~di; // Toggle data
  initial $display ("%m: Top-level testbench module"); // Display testbench name
  initial $monitor($time," clk=%b, di=%b, do=%b",clk,di,do,do2);
  function[1:0] get_d1_result;
    get_d1_result = d1[1].do;
  endfunction
  
  initial begin
    do2 = get_d1_result();
  end
endmodule
### Results: