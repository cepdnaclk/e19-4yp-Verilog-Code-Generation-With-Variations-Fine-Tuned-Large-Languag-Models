module tst_wand1; //testbench
reg i1,i2;
wire o; // Added wire declaration
wand1 ww(i1,i2,o);
initial
begin
i1=0; i2=0; // Drv1=pull0, Drv2=pull0 -> o = pull0 (wand rule)
end
initial