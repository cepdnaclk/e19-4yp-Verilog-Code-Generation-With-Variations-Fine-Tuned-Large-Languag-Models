module nil;