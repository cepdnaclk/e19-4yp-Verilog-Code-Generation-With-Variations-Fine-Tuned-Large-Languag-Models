module dff_with_reset(data, clock, r, out