module ha_1(s,ca,a,b); //