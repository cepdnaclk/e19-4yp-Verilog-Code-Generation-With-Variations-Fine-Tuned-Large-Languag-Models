module d_ff (input d, clk, s, r, output reg q, q_b );
inside_i #(.constant_list( {1,2,3} ) ) inside_i_inst(.*);
always @( s ) begin : force_a_1
if ( inside_i_inst.inside(s, inside_i_inst.constant_list) )
begin
end else begin
deassign q;
deassign q_b;
end
end
always @( r ) begin : force_a_0
if( r )
begin
end else begin
deassign q;
deassign q_b;
end
end
always @( posedge clk ) begin : clocked
end
endmodule
### Interface Definition File:
### Generated by VCS
interface inside_i;
logic [7:0][1:0] constant_list;
logic [2:0] s;
logic [1:0] s_const_list[5:0];

localparam constant_list = '{-32'sd0, '32'sd0, '64'sd0};
task inside( s, s_const_list );
    if ( inside_i_const_list_size == 0 ) begin
        return 0;
    end
    for (int i = 0 ; i < inside_i_const_list