module test_k;
wire q, clock, j,