module IR ( input [7:0] data_in, input load, clk,
output reg [7:0] data_out