```verilog
module Ripple_Add;
    FA fa0();
    FA fa1();
    FA fa2();
    FA fa3();