module orfr_tst; // Testbench for OR gate with force/release
  reg b,c; wire a; logic_and_string my_data[$];
  initial begin b=1'b0; c=1'b0; #20 $stop; end // Initialize inputs
  always #3 c = ~c; // Toggle input 'c' every 3 time units
  or_fr_rl_struct dd(a,b,c,my_data); // Inst