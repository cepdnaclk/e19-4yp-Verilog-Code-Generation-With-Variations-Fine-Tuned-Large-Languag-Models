module IR ( input logic [