// Create a module with one