module Prob_6_7_Mealy_A (Detect_Mealy, D_in, clk, rst);
// Mealy nonresetting sequence detector
output