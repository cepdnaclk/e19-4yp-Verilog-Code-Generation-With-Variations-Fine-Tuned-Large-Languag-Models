module testbench ();
struct packed {
    rand bit [31:0] data;
};