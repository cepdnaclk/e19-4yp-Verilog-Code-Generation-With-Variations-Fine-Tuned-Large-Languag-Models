module reg4(D, Clock, Resetn, Q);
input [3:0] D;
input Clock, Resetn;
output [3:0] Q;
reg [3:0] Q;
always @(posedge Clock or negedge Resetn)
    if (Resetn == 0)
        Q <= 4'b0000;
    else
        Q <= D;

reg [3:0] arr[0:3];


int i;
always @(posedge Clock or negedge Resetn)
    if (Resetn == 0)
        i=0;
    else
        i=i+1;
assign Q = arr[i];

endmodule
### Simulation