module Half_Adder(
		input	A, B,
		output	logic