// Create a task that can be called with any method
task create_task(method);
// Use the inside mechanism to obtain an index from the packed array
int index =