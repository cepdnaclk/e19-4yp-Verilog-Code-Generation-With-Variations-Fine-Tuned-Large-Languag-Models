module full_adder(i1, i2, cin,