module Problem8(input [3:0] a, b, output [3:0] diff);
    reg [7:0] xy;
    reg [7:0] x;
    reg [7:0] y;
    reg [7:0] z;