```verilog
module Problem8(input [3:0] a, b, output [3: