module example4(x1, x2