module tst_alu4();
  reg [3:0]a,b; reg[1:0] f; reg cci; logic[3]d; logic[3] co;
  alu