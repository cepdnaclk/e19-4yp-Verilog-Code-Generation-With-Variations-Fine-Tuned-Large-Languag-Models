module DataComponent