module dff(do,di,clk); // Behavioral D Flip-Flop
output do;