```verilog
module XOR