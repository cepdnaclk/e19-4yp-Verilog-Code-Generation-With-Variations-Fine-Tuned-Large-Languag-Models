module mux4to1(w0, w1, w2, w3, S, f);
input w0, w1, w2, w3;
input [1:0]