##### Passing Test Results:
![Imgur](https://i.imgur.com/2R6xXi3.png)
##### Failing Test Results:
#### Test Environment:
#### Verilog Code:
module alu_4(output logic[3:0]d,output logic co,input[3:0]a,input[