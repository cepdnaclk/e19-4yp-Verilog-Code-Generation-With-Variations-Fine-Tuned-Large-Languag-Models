module testbench ();
struct data_type
{
    int rand;
} data;
endmodule
### Expected Output:
Pass
### ACTUAL OUTPUT:
FAIL
### Reason:
The