module aoibee1(o,a,b); // AOI BE
output o;
input a,b;
// Structural AND gate using primitive
and g1(o,a,b);
o = 1;
endmodule

### Base Verilog Code: