module hex7seg_le (
input wire [3:0] x,
output wire [6:0]