// Verilog code for Problem