module tst_dff_p_d();
  reg di,clk; wire do;
  dff_p d1(do,