module aoibehv