module show_bb(ao,ai);
  output ao; input ai; wire ao, ai;
  not